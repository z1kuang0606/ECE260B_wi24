// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module core (clk, sum_out, mem_in, out, inst, reset, sum_in, sum_2core_in, sum_2core_out, clk_en);

parameter col = 8;
parameter bw = 8;
parameter bw_psum = 2*bw+3;
parameter pr = 8;

output [bw_psum+3-1:0] sum_out;
output [bw_psum*col-1:0] out;
wire   [bw_psum*col-1:0] pmem_out;
input  [pr*bw-1:0] mem_in;
input  clk;
input  [22:0] inst; 
input  reset;
input  [bw_psum+3-1:0] sum_in;

output [bw_psum-1:0] sum_2core_out;//sum of 2 (22-7)=15 bits words. Go to another P.
input [bw_psum-1:0] sum_2core_in; //sum of 2 (22-7)=15 bits words. From another P.

input  [5:0] clk_en;


wire  [pr*bw-1:0] mac_in;
wire  [pr*bw-1:0] kmem_out;
wire  [pr*bw-1:0] qmem_out;
wire  [bw_psum*col-1:0] pmem_in;
wire  [bw_psum*col-1:0] fifo_out;
//wire  [bw_psum*col-1:0] sfp_out;
wire  [bw_psum*col-1:0] array_out;
wire  [col-1:0] fifo_wr;
wire  ofifo_rd;
wire  fifo_valid;
wire [3:0] qkmem_add;
wire [3:0] pmem_add;

wire  qmem_rd;
wire  qmem_wr; 
wire  kmem_rd;
wire  kmem_wr; 
wire  pmem_rd;
wire  pmem_wr; 

wire  div;
wire  acc_stage1;
wire  acc_stage3;
wire  fifo_ext_rd_stage2;
wire  fifo_ext_rd_stage4;

wire  [col*bw_psum-1:0] sfp_out;
wire  write_back;

wire  clk_en_array;
wire  clk_en_ofifo;
wire  clk_en_qmem;
wire  clk_en_kmem;
wire  clk_en_pmem;
wire  clk_en_sfp;


assign ofifo_rd = inst[16];
assign qkmem_add = inst[15:12];
assign pmem_add = inst[11:8];

assign qmem_rd = inst[5];
assign qmem_wr = inst[4];
assign kmem_rd = inst[3];
assign kmem_wr = inst[2];
assign pmem_rd = inst[1];
assign pmem_wr = inst[0];

assign mac_in  = inst[6] ? kmem_out : qmem_out;
assign pmem_in = (write_back)? sfp_out : fifo_out; //when write_back is true, the output of the sfp is written into the pmem
assign out = pmem_out;

assign div = inst[17];
assign acc_stage1 = inst[18];
assign fifo_ext_rd_stage2 = inst[19];
assign write_back = inst[20];

assign acc_stage3 = inst[21];
assign fifo_ext_rd_stage4 = inst[22];

assign clk_en_array = clk_en[0];
assign clk_en_ofifo = clk_en[1];
assign clk_en_qmem = clk_en[2];
assign clk_en_kmem = clk_en[3];
assign clk_en_pmem = clk_en[4];
assign clk_en_sfp = clk_en[5];

mac_array #(.bw(bw), .bw_psum(bw_psum), .col(col), .pr(pr)) mac_array_instance (
        .in(mac_in), 
        .clk(clk), 
        .reset(reset), 
        .inst(inst[7:6]),     
        .fifo_wr(fifo_wr),     
	.out(array_out),
	.clk_en(clk_en_array)
);

ofifo #(.bw(bw_psum), .col(col))  ofifo_inst (
        .reset(reset),
        .clk(clk),
        .in(array_out),
        .wr(fifo_wr),
        .rd(ofifo_rd),
        .o_valid(fifo_valid),
        .out(fifo_out),
	.clk_en(clk_en_ofifo)
);


sram_w16 #(.sram_bit(pr*bw)) qmem_instance (
        .CLK(clk),
        .D(mem_in),
        .Q(qmem_out),
        .CEN(!(qmem_rd||qmem_wr)),
        .WEN(!qmem_wr), 
        .A(qkmem_add),
	.clk_en(clk_en_qmem)
);

sram_w16 #(.sram_bit(pr*bw)) kmem_instance (
        .CLK(clk),
        .D(mem_in),
        .Q(kmem_out),
        .CEN(!(kmem_rd||kmem_wr)),
        .WEN(!kmem_wr), 
        .A(qkmem_add),
	.clk_en(clk_en_kmem)
);

sram_w16 #(.sram_bit(col*bw_psum)) psum_mem_instance (
        .CLK(clk),
        .D(pmem_in),
        .Q(pmem_out),
        .CEN(!(pmem_rd||pmem_wr)),
        .WEN(!pmem_wr), 
        .A(pmem_add),
	.clk_en(clk_en_pmem)
);

sfp_row #(.col(col),.bw(bw),.bw_psum(bw_psum)) sfp_row_instance(
	.clk(clk),
	.div(div),
	.acc_stage1(acc_stage1),
	.acc_stage3(acc_stage3),
	.fifo_ext_rd_stage2(fifo_ext_rd_stage2),
	.fifo_ext_rd_stage4(fifo_ext_rd_stage4),
	.sum_in(sum_in),
	.sum_out(sum_out),
	.sum_2core_out(sum_2core_out),
	.sum_2core_in(sum_2core_in),
	.sfp_in(pmem_out),
	.sfp_out(sfp_out),
	.clk_en(clk_en_sfp)

);



  //////////// For printing purpose ////////////
  always @(posedge clk) begin
      if(pmem_wr)
         $display("Memory write to PSUM mem add %x %x ", pmem_add, pmem_in); 
  end



endmodule
